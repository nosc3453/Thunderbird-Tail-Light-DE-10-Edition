parameter IDLE = 1;
parameter HAZARD = 2;
parameter RIGHT = 3;
parameter LEFT = 4;